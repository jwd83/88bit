/*

The ShinyRock16

My ISA Defined here:

https://docs.google.com/spreadsheets/d/e/2PACX-1vTi-MPLhr4D1eNBMzdLoQ9VZIzOb1GxG1HfwbSVVtuh3BAOuYNPyyuVTR7AJ4V3hfcSsUTbSlYO6jC3/pubhtml

*/