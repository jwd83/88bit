// a collection of 8 bit adders and their components

// half adder
// full adder
// 4 bit ripple carry adder
// 8 bit ripple carry adder
// 8 bit carry select adder, zoom, zoom
