/*

The ShinyRock16

*/